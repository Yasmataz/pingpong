--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   00:05:23 12/05/2020
-- Design Name:   
-- Module Name:   C:/Users/Yasamin/Documents/Classes/COE758/Spartan3E-master/refresh_test.vhd
-- Project Name:  VGA
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: refreshClk
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY refresh_test IS
END refresh_test;
 
ARCHITECTURE behavior OF refresh_test IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT refreshClk
    PORT(
         clk : IN  std_logic;
         p_clk : IN  std_logic;
         rcount : OUT  integer;
         rclk : OUT  std_logic
        );
    END COMPONENT;
    

   --Inputs
   signal clk : std_logic := '0';
   signal p_clk : std_logic := '0';

 	--Outputs
   signal rcount : integer;
   signal rclk : std_logic;

   -- Clock period definitions
   constant clk_period : time := 10 ns;
   constant p_clk_period : time := 20 ns;
   constant rclk_period : time := 10 ns;
 
BEGIN
  
	-- Instantiate the Unit Under Test (UUT)
   uut: refreshClk PORT MAP (
          clk => clk,
          p_clk => p_clk,
          rcount => rcount,
          rclk => rclk
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 
   p_clk_process :process
   begin
		p_clk <= '0';
		wait for p_clk_period/2;
		p_clk <= '1';
		wait for p_clk_period/2;
   end process;
 
   rclk_process :process
   begin
		rclk <= '0';
		wait for rclk_period/2;
		rclk <= '1';
		wait for rclk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	

      wait for clk_period*10;

      -- insert stimulus here 

      wait;
   end process;

END;
